// CPU1_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU1_tb (
	);

	wire        cpu1_inst_clk_bfm_clk_clk; // CPU1_inst_clk_bfm:clk -> CPU1_inst:clk_clk
	wire  [1:0] cpu1_inst_leds_export;     // CPU1_inst:leds_export -> CPU1_inst_leds_bfm:sig_export

	CPU1 cpu1_inst (
		.clk_clk     (cpu1_inst_clk_bfm_clk_clk), //  clk.clk
		.leds_export (cpu1_inst_leds_export)      // leds.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) cpu1_inst_clk_bfm (
		.clk (cpu1_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm cpu1_inst_leds_bfm (
		.sig_export (cpu1_inst_leds_export)  // conduit.export
	);

endmodule
