
module unsaved (
	onchip_memory2_0_clk1_clk);	

	input		onchip_memory2_0_clk1_clk;
endmodule
