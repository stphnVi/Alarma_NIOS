// CPU1.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU1 (
		output wire       buz_export,          //          buz.export
		input  wire       clk_clk,             //          clk.clk
		input  wire       hours_export,        //        hours.export
		output wire [1:0] leds_export,         //         leds.export
		input  wire       minutes_export,      //      minutes.export
		input  wire       off_export,          //          off.export
		input  wire       reset_reset_n,       //        reset.reset_n
		output wire [6:0] s1_export,           //           s1.export
		output wire [6:0] s2_export,           //           s2.export
		output wire [6:0] s3_export,           //           s3.export
		output wire [6:0] s4_export,           //           s4.export
		input  wire       set_alarm_export,    //    set_alarm.export
		input  wire       set_clock_export,    //    set_clock.export
		input  wire       switch_reset_export  // switch_reset.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [13:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [13:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_pio_leds_0_s1_chipselect;                  // mm_interconnect_0:pio_leds_0_s1_chipselect -> pio_leds_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_leds_0_s1_readdata;                    // pio_leds_0:readdata -> mm_interconnect_0:pio_leds_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_leds_0_s1_address;                     // mm_interconnect_0:pio_leds_0_s1_address -> pio_leds_0:address
	wire         mm_interconnect_0_pio_leds_0_s1_write;                       // mm_interconnect_0:pio_leds_0_s1_write -> pio_leds_0:write_n
	wire  [31:0] mm_interconnect_0_pio_leds_0_s1_writedata;                   // mm_interconnect_0:pio_leds_0_s1_writedata -> pio_leds_0:writedata
	wire         mm_interconnect_0_pio_s4_s1_chipselect;                      // mm_interconnect_0:pio_s4_s1_chipselect -> pio_s4:chipselect
	wire  [31:0] mm_interconnect_0_pio_s4_s1_readdata;                        // pio_s4:readdata -> mm_interconnect_0:pio_s4_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_s4_s1_address;                         // mm_interconnect_0:pio_s4_s1_address -> pio_s4:address
	wire         mm_interconnect_0_pio_s4_s1_write;                           // mm_interconnect_0:pio_s4_s1_write -> pio_s4:write_n
	wire  [31:0] mm_interconnect_0_pio_s4_s1_writedata;                       // mm_interconnect_0:pio_s4_s1_writedata -> pio_s4:writedata
	wire         mm_interconnect_0_pio_s1_s1_chipselect;                      // mm_interconnect_0:pio_s1_s1_chipselect -> pio_s1:chipselect
	wire  [31:0] mm_interconnect_0_pio_s1_s1_readdata;                        // pio_s1:readdata -> mm_interconnect_0:pio_s1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_s1_s1_address;                         // mm_interconnect_0:pio_s1_s1_address -> pio_s1:address
	wire         mm_interconnect_0_pio_s1_s1_write;                           // mm_interconnect_0:pio_s1_s1_write -> pio_s1:write_n
	wire  [31:0] mm_interconnect_0_pio_s1_s1_writedata;                       // mm_interconnect_0:pio_s1_s1_writedata -> pio_s1:writedata
	wire         mm_interconnect_0_pio_s2_s1_chipselect;                      // mm_interconnect_0:pio_s2_s1_chipselect -> pio_s2:chipselect
	wire  [31:0] mm_interconnect_0_pio_s2_s1_readdata;                        // pio_s2:readdata -> mm_interconnect_0:pio_s2_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_s2_s1_address;                         // mm_interconnect_0:pio_s2_s1_address -> pio_s2:address
	wire         mm_interconnect_0_pio_s2_s1_write;                           // mm_interconnect_0:pio_s2_s1_write -> pio_s2:write_n
	wire  [31:0] mm_interconnect_0_pio_s2_s1_writedata;                       // mm_interconnect_0:pio_s2_s1_writedata -> pio_s2:writedata
	wire         mm_interconnect_0_pio_s3_s1_chipselect;                      // mm_interconnect_0:pio_s3_s1_chipselect -> pio_s3:chipselect
	wire  [31:0] mm_interconnect_0_pio_s3_s1_readdata;                        // pio_s3:readdata -> mm_interconnect_0:pio_s3_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_s3_s1_address;                         // mm_interconnect_0:pio_s3_s1_address -> pio_s3:address
	wire         mm_interconnect_0_pio_s3_s1_write;                           // mm_interconnect_0:pio_s3_s1_write -> pio_s3:write_n
	wire  [31:0] mm_interconnect_0_pio_s3_s1_writedata;                       // mm_interconnect_0:pio_s3_s1_writedata -> pio_s3:writedata
	wire         mm_interconnect_0_pio_buzz_0_s1_chipselect;                  // mm_interconnect_0:pio_buzz_0_s1_chipselect -> pio_buzz_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_buzz_0_s1_readdata;                    // pio_buzz_0:readdata -> mm_interconnect_0:pio_buzz_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_buzz_0_s1_address;                     // mm_interconnect_0:pio_buzz_0_s1_address -> pio_buzz_0:address
	wire         mm_interconnect_0_pio_buzz_0_s1_write;                       // mm_interconnect_0:pio_buzz_0_s1_write -> pio_buzz_0:write_n
	wire  [31:0] mm_interconnect_0_pio_buzz_0_s1_writedata;                   // mm_interconnect_0:pio_buzz_0_s1_writedata -> pio_buzz_0:writedata
	wire  [31:0] mm_interconnect_0_pio_switch_off_s1_readdata;                // pio_switch_off:readdata -> mm_interconnect_0:pio_switch_off_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_switch_off_s1_address;                 // mm_interconnect_0:pio_switch_off_s1_address -> pio_switch_off:address
	wire  [31:0] mm_interconnect_0_pio_set_alarm_s1_readdata;                 // pio_set_alarm:readdata -> mm_interconnect_0:pio_set_alarm_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_set_alarm_s1_address;                  // mm_interconnect_0:pio_set_alarm_s1_address -> pio_set_alarm:address
	wire  [31:0] mm_interconnect_0_pio_switch_clock_s1_readdata;              // pio_switch_clock:readdata -> mm_interconnect_0:pio_switch_clock_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_switch_clock_s1_address;               // mm_interconnect_0:pio_switch_clock_s1_address -> pio_switch_clock:address
	wire  [31:0] mm_interconnect_0_pio_switch_reset_s1_readdata;              // pio_switch_reset:readdata -> mm_interconnect_0:pio_switch_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_switch_reset_s1_address;               // mm_interconnect_0:pio_switch_reset_s1_address -> pio_switch_reset:address
	wire         mm_interconnect_0_pio_button_hours_s1_chipselect;            // mm_interconnect_0:pio_button_hours_s1_chipselect -> pio_button_hours:chipselect
	wire  [31:0] mm_interconnect_0_pio_button_hours_s1_readdata;              // pio_button_hours:readdata -> mm_interconnect_0:pio_button_hours_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_button_hours_s1_address;               // mm_interconnect_0:pio_button_hours_s1_address -> pio_button_hours:address
	wire         mm_interconnect_0_pio_button_hours_s1_write;                 // mm_interconnect_0:pio_button_hours_s1_write -> pio_button_hours:write_n
	wire  [31:0] mm_interconnect_0_pio_button_hours_s1_writedata;             // mm_interconnect_0:pio_button_hours_s1_writedata -> pio_button_hours:writedata
	wire         mm_interconnect_0_pio_button_minutes_s1_chipselect;          // mm_interconnect_0:pio_button_minutes_s1_chipselect -> pio_button_minutes:chipselect
	wire  [31:0] mm_interconnect_0_pio_button_minutes_s1_readdata;            // pio_button_minutes:readdata -> mm_interconnect_0:pio_button_minutes_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_button_minutes_s1_address;             // mm_interconnect_0:pio_button_minutes_s1_address -> pio_button_minutes:address
	wire         mm_interconnect_0_pio_button_minutes_s1_write;               // mm_interconnect_0:pio_button_minutes_s1_write -> pio_button_minutes:write_n
	wire  [31:0] mm_interconnect_0_pio_button_minutes_s1_writedata;           // mm_interconnect_0:pio_button_minutes_s1_writedata -> pio_button_minutes:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // pio_button_hours:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // pio_button_minutes:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // timer_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, pio_button_hours:reset_n, pio_button_minutes:reset_n, pio_buzz_0:reset_n, pio_leds_0:reset_n, pio_s1:reset_n, pio_s2:reset_n, pio_s3:reset_n, pio_s4:reset_n, pio_set_alarm:reset_n, pio_switch_clock:reset_n, pio_switch_off:reset_n, pio_switch_reset:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]

	CPU1_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	CPU1_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	CPU1_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	CPU1_pio_button_hours pio_button_hours (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_pio_button_hours_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_button_hours_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_button_hours_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_button_hours_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_button_hours_s1_readdata),   //                    .readdata
		.in_port    (hours_export),                                     // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                          //                 irq.irq
	);

	CPU1_pio_button_hours pio_button_minutes (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_button_minutes_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_button_minutes_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_button_minutes_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_button_minutes_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_button_minutes_s1_readdata),   //                    .readdata
		.in_port    (minutes_export),                                     // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                            //                 irq.irq
	);

	CPU1_pio_buzz_0 pio_buzz_0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_buzz_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_buzz_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_buzz_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_buzz_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_buzz_0_s1_readdata),   //                    .readdata
		.out_port   (buz_export)                                  // external_connection.export
	);

	CPU1_pio_leds_0 pio_leds_0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_leds_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_leds_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_leds_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_leds_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_leds_0_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                                 // external_connection.export
	);

	CPU1_pio_s1 pio_s1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_pio_s1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_s1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_s1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_s1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_s1_s1_readdata),   //                    .readdata
		.out_port   (s1_export)                               // external_connection.export
	);

	CPU1_pio_s1 pio_s2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_pio_s2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_s2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_s2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_s2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_s2_s1_readdata),   //                    .readdata
		.out_port   (s2_export)                               // external_connection.export
	);

	CPU1_pio_s1 pio_s3 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_pio_s3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_s3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_s3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_s3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_s3_s1_readdata),   //                    .readdata
		.out_port   (s3_export)                               // external_connection.export
	);

	CPU1_pio_s1 pio_s4 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_pio_s4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_s4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_s4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_s4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_s4_s1_readdata),   //                    .readdata
		.out_port   (s4_export)                               // external_connection.export
	);

	CPU1_pio_set_alarm pio_set_alarm (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_pio_set_alarm_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_set_alarm_s1_readdata), //                    .readdata
		.in_port  (set_alarm_export)                             // external_connection.export
	);

	CPU1_pio_set_alarm pio_switch_clock (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_pio_switch_clock_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_switch_clock_s1_readdata), //                    .readdata
		.in_port  (set_clock_export)                                // external_connection.export
	);

	CPU1_pio_set_alarm pio_switch_off (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pio_switch_off_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_switch_off_s1_readdata), //                    .readdata
		.in_port  (off_export)                                    // external_connection.export
	);

	CPU1_pio_set_alarm pio_switch_reset (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_pio_switch_reset_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_switch_reset_s1_readdata), //                    .readdata
		.in_port  (switch_reset_export)                             // external_connection.export
	);

	CPU1_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	CPU1_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                              //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.pio_button_hours_s1_address                    (mm_interconnect_0_pio_button_hours_s1_address),               //                      pio_button_hours_s1.address
		.pio_button_hours_s1_write                      (mm_interconnect_0_pio_button_hours_s1_write),                 //                                         .write
		.pio_button_hours_s1_readdata                   (mm_interconnect_0_pio_button_hours_s1_readdata),              //                                         .readdata
		.pio_button_hours_s1_writedata                  (mm_interconnect_0_pio_button_hours_s1_writedata),             //                                         .writedata
		.pio_button_hours_s1_chipselect                 (mm_interconnect_0_pio_button_hours_s1_chipselect),            //                                         .chipselect
		.pio_button_minutes_s1_address                  (mm_interconnect_0_pio_button_minutes_s1_address),             //                    pio_button_minutes_s1.address
		.pio_button_minutes_s1_write                    (mm_interconnect_0_pio_button_minutes_s1_write),               //                                         .write
		.pio_button_minutes_s1_readdata                 (mm_interconnect_0_pio_button_minutes_s1_readdata),            //                                         .readdata
		.pio_button_minutes_s1_writedata                (mm_interconnect_0_pio_button_minutes_s1_writedata),           //                                         .writedata
		.pio_button_minutes_s1_chipselect               (mm_interconnect_0_pio_button_minutes_s1_chipselect),          //                                         .chipselect
		.pio_buzz_0_s1_address                          (mm_interconnect_0_pio_buzz_0_s1_address),                     //                            pio_buzz_0_s1.address
		.pio_buzz_0_s1_write                            (mm_interconnect_0_pio_buzz_0_s1_write),                       //                                         .write
		.pio_buzz_0_s1_readdata                         (mm_interconnect_0_pio_buzz_0_s1_readdata),                    //                                         .readdata
		.pio_buzz_0_s1_writedata                        (mm_interconnect_0_pio_buzz_0_s1_writedata),                   //                                         .writedata
		.pio_buzz_0_s1_chipselect                       (mm_interconnect_0_pio_buzz_0_s1_chipselect),                  //                                         .chipselect
		.pio_leds_0_s1_address                          (mm_interconnect_0_pio_leds_0_s1_address),                     //                            pio_leds_0_s1.address
		.pio_leds_0_s1_write                            (mm_interconnect_0_pio_leds_0_s1_write),                       //                                         .write
		.pio_leds_0_s1_readdata                         (mm_interconnect_0_pio_leds_0_s1_readdata),                    //                                         .readdata
		.pio_leds_0_s1_writedata                        (mm_interconnect_0_pio_leds_0_s1_writedata),                   //                                         .writedata
		.pio_leds_0_s1_chipselect                       (mm_interconnect_0_pio_leds_0_s1_chipselect),                  //                                         .chipselect
		.pio_s1_s1_address                              (mm_interconnect_0_pio_s1_s1_address),                         //                                pio_s1_s1.address
		.pio_s1_s1_write                                (mm_interconnect_0_pio_s1_s1_write),                           //                                         .write
		.pio_s1_s1_readdata                             (mm_interconnect_0_pio_s1_s1_readdata),                        //                                         .readdata
		.pio_s1_s1_writedata                            (mm_interconnect_0_pio_s1_s1_writedata),                       //                                         .writedata
		.pio_s1_s1_chipselect                           (mm_interconnect_0_pio_s1_s1_chipselect),                      //                                         .chipselect
		.pio_s2_s1_address                              (mm_interconnect_0_pio_s2_s1_address),                         //                                pio_s2_s1.address
		.pio_s2_s1_write                                (mm_interconnect_0_pio_s2_s1_write),                           //                                         .write
		.pio_s2_s1_readdata                             (mm_interconnect_0_pio_s2_s1_readdata),                        //                                         .readdata
		.pio_s2_s1_writedata                            (mm_interconnect_0_pio_s2_s1_writedata),                       //                                         .writedata
		.pio_s2_s1_chipselect                           (mm_interconnect_0_pio_s2_s1_chipselect),                      //                                         .chipselect
		.pio_s3_s1_address                              (mm_interconnect_0_pio_s3_s1_address),                         //                                pio_s3_s1.address
		.pio_s3_s1_write                                (mm_interconnect_0_pio_s3_s1_write),                           //                                         .write
		.pio_s3_s1_readdata                             (mm_interconnect_0_pio_s3_s1_readdata),                        //                                         .readdata
		.pio_s3_s1_writedata                            (mm_interconnect_0_pio_s3_s1_writedata),                       //                                         .writedata
		.pio_s3_s1_chipselect                           (mm_interconnect_0_pio_s3_s1_chipselect),                      //                                         .chipselect
		.pio_s4_s1_address                              (mm_interconnect_0_pio_s4_s1_address),                         //                                pio_s4_s1.address
		.pio_s4_s1_write                                (mm_interconnect_0_pio_s4_s1_write),                           //                                         .write
		.pio_s4_s1_readdata                             (mm_interconnect_0_pio_s4_s1_readdata),                        //                                         .readdata
		.pio_s4_s1_writedata                            (mm_interconnect_0_pio_s4_s1_writedata),                       //                                         .writedata
		.pio_s4_s1_chipselect                           (mm_interconnect_0_pio_s4_s1_chipselect),                      //                                         .chipselect
		.pio_set_alarm_s1_address                       (mm_interconnect_0_pio_set_alarm_s1_address),                  //                         pio_set_alarm_s1.address
		.pio_set_alarm_s1_readdata                      (mm_interconnect_0_pio_set_alarm_s1_readdata),                 //                                         .readdata
		.pio_switch_clock_s1_address                    (mm_interconnect_0_pio_switch_clock_s1_address),               //                      pio_switch_clock_s1.address
		.pio_switch_clock_s1_readdata                   (mm_interconnect_0_pio_switch_clock_s1_readdata),              //                                         .readdata
		.pio_switch_off_s1_address                      (mm_interconnect_0_pio_switch_off_s1_address),                 //                        pio_switch_off_s1.address
		.pio_switch_off_s1_readdata                     (mm_interconnect_0_pio_switch_off_s1_readdata),                //                                         .readdata
		.pio_switch_reset_s1_address                    (mm_interconnect_0_pio_switch_reset_s1_address),               //                      pio_switch_reset_s1.address
		.pio_switch_reset_s1_readdata                   (mm_interconnect_0_pio_switch_reset_s1_readdata),              //                                         .readdata
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect)                      //                                         .chipselect
	);

	CPU1_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
